

module not32(OUT, IN);

input [31:0] IN;
output [31:0] OUT;

not not0(OUT[0], IN[0]);
not not1(OUT[1], IN[1]);
not not2(OUT[2], IN[2]);
not not3(OUT[3], IN[3]);
not not4(OUT[4], IN[4]);
not not5(OUT[5], IN[5]);
not not6(OUT[6], IN[6]);
not not7(OUT[7], IN[7]);
not not8(OUT[8], IN[8]);
not not9(OUT[9], IN[9]);
not not10(OUT[10], IN[10]);
not not11(OUT[11], IN[11]);
not not12(OUT[12], IN[12]);
not not13(OUT[13], IN[13]);
not not14(OUT[14], IN[14]);
not not15(OUT[15], IN[15]);
not not16(OUT[16], IN[16]);
not not17(OUT[17], IN[17]);
not not18(OUT[18], IN[18]);
not not19(OUT[19], IN[19]);
not not20(OUT[20], IN[20]);
not not21(OUT[21], IN[21]);
not not22(OUT[22], IN[22]);
not not23(OUT[23], IN[23]);
not not24(OUT[24], IN[24]);
not not25(OUT[25], IN[25]);
not not26(OUT[26], IN[26]);
not not27(OUT[27], IN[27]);
not not28(OUT[28], IN[28]);
not not29(OUT[29], IN[29]);
not not30(OUT[30], IN[30]);
not not31(OUT[31], IN[31]);

endmodule